***y = (A+(B+C).D+E)'	***
VD 10 0 dc 2.5V
VGA 1 0 pulse (5 0 0 0 0 2.5 5)
VGB 2 0 pulse (7.5 0 0 0 0 5 10)
VGC 3 0 pulse (10 0 0 0 0 7.5 15)
VGD 4 0 pulse (12.5 0 0 0 0 10 20)
VGE 5 0 pulse (15 0 0 0 0 12.5 25)

.model nmod nmos level=54 version=4.7
M1 7 1 0 0 nmod w=10u l=1u
M2 6 2 0 0 nmod w=10u l=1u
M3 6 3 0 0 nmod w=10u l=1u
M4 7 4 6 6 nmod w=10u l=1u
M5 7 5 0 0 nmod w=10u l=1u

.model pmod pmos level=54 version=4.7
M6 8 1 9 9 pmod w=10u l=1u
M7 9 2 11 11 pmod w=10u l=1u
M8 11 3 10 10 pmod w=10u l=1u
M9 9 4 10 10 pmod w=10u l=1u
M10 7 5 8 8 pmod w=10u l=1u

.tran 0.1 80
.control
run
plot V(4) V(1) V(2) V(3) V(5) V(7) 
.endc
.end

