*** Transmission Gate***

.subckt cmos_inv 1 2 3
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 3 1 0 0 nmod w=100u l=10u
M2 3 1 2 2 pmod w=100u l=10u
.ends

.subckt cmos_tran 1 2 3 4
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 1 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 pmod w=100u l=10u
.ends

VA 10 0 pulse(5 0 0 0 0 10 20)
VB 11 0 dc 5V
Vdd 2 0 dc 10V

xa 10 2 12 cmos_inv
xb 11 2 13 cmos_inv

xab_bar 12 11 13 14 cmos_tran
xa_barb 10 13 11 14 cmos_tran

.tran 0.1 100 
.control
run
plot V(10) V(14) V(12)
.endc
.end