***y = a.b.c+d(Pass Transistor Technique)***
.subckt pass_or 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 1 3 4 4 nmod w=100u l=10u
M2 2 2 4 4 nmod w=100u l=10u
.ends

.subckt pass_and 1 2 3 4
.model nmod nmos level=54 version=4.7
M1 1 2 4 4 nmod w=100u l=10u
M2 2 3 4 4 nmod w=100u l=10u
.ends

.subckt cmos_inv 1 2 3
.model nmod nmos level=54 version=4.7
.model pmod pmos level=54 version=4.7
M1 3 1 0 0 nmod w=100u l=10u
M2 3 1 2 2 pmod w=100u l=10u
.ends

VA 10 0 pulse(5 0 0 0 0 10 20)
VB 11 0 pulse(10 0 0 0 0 15 25)
VC 12 0 pulse(15 0 0 0 0 20 30)
VD 13 0 dc 0V
Vdd 2 0 dc 5V

xa 10 2 14 cmos_inv
xc 12 2 15 cmos_inv
xd 13 2 16 cmos_inv

xaandb 11 10 14 17 pass_and
xabandc 17 12 15 18 pass_and
xabcord 18 13 16 19 pass_or

.tran 0.1 200 
.control
run
plot V(10) V(19) V(11) V(12)
.endc
.end