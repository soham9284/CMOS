***2 input NAND Gate***
VGA 3 0 pulse (7.5 0 0 0 0 5 10)
VGB 1 0 pulse (10 0 0 0 0 10 20)
VD 5 0 dc 5V

.model nmod nmos level=54 version=4.7
M1 2 1 0 0 nmod w=10u l=1u
M2 4 3 2 2 nmod w=10u l=1u

.model pmod pmos level=54 version=4.7
M3 4 1 5 5 pmod w=10u l=1u
M4 4 3 5 5 pmod w=10u l=1u

.tran 0.1 40

.control
run
plot V(4) V(3) V(1)
.endc
.end
