***COMMON SOURCE AMPLIFIER***
VDD 2 0 dc 1.2V
VB 4 0 dc 0.6V
VIN 5 0 SIN (0.6 0.1 200M)

.model nmod nmos level=54 version=4.7
M1 1 4 0 0 nmod w=5u l=0.1u
M2 3 5 0 0 nmod w=5u l=0.1u

.model pmod pmos level=54 version=4.7
M3 2 1 1 1 pmod w=5u l=0.1u
M4 2 1 3 3 pmod w=5u l=0.1u

.tran 0.1 80
.control
run
plot V(5) V(3)  
.endc
.end
